.circuit
I1   1 GND  dc 3
R1   2   1  6
R2   2 GND  9
.end
